magic
tech sky130A
magscale 1 2
timestamp 1624128865
<< metal2 >>
rect 466000 700695 469800 700700
rect 393100 697295 417800 697300
rect 120800 694095 360500 694100
rect 120796 690305 120805 694095
rect 124595 690305 360500 694095
rect 120800 690300 360500 690305
rect 68805 677000 72395 677004
rect 68800 676995 350600 677000
rect 68800 673405 68805 676995
rect 72395 673405 350600 676995
rect 68800 673400 350600 673405
rect 68805 673396 72395 673400
rect 16807 662188 340793 662193
rect 16803 658612 16812 662188
rect 20388 658612 340793 662188
rect 16807 658607 340793 658612
rect 337207 653407 340793 658607
rect 299570 644548 328604 644593
rect 299570 644520 329043 644548
rect 299570 644481 328604 644520
rect -2 1 1 610629
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 644481
rect 339127 643400 339927 653407
rect 347000 653200 350600 673400
rect 349117 643600 349917 653200
rect 356700 653100 360500 690300
rect 393100 693505 414005 697295
rect 417795 693505 417804 697295
rect 465996 696905 466005 700695
rect 469795 696905 469804 700695
rect 393100 693500 417800 693505
rect 359107 642400 359907 653100
rect 393100 652500 396900 693500
rect 466000 689700 469800 696905
rect 406900 685900 469800 689700
rect 554703 691292 570997 691297
rect 554703 687508 567208 691292
rect 570992 687508 571001 691292
rect 554703 687503 570997 687508
rect 406900 652500 410700 685900
rect 554703 682097 558497 687503
rect 573705 682600 577895 682604
rect 418000 678303 558497 682097
rect 564100 682595 577900 682600
rect 564100 678405 573705 682595
rect 577895 678405 577900 682595
rect 564100 678400 577900 678405
rect 418000 652703 421497 678303
rect 564100 672700 568300 678400
rect 573705 678396 577895 678400
rect 426300 668500 568300 672700
rect 394109 642800 394909 652500
rect 409131 642400 409931 652500
rect 418921 642600 420121 652703
rect 426300 652700 430500 668500
rect 427875 642600 429075 652700
rect 509944 644548 510056 644589
rect 509440 644520 510056 644548
rect 509944 644256 510056 644520
rect 509944 644144 576270 644256
rect 510001 637291 572724 637403
rect 510001 637252 510113 637291
rect 509440 637224 510113 637252
rect 510001 637193 510113 637224
rect 303116 634468 328609 634495
rect 303116 634440 329033 634468
rect 303116 634383 328609 634440
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 634383
rect 510002 629956 510114 629998
rect 509399 629928 510114 629956
rect 510002 629431 510114 629928
rect 510002 629319 569178 629431
rect 306662 624484 328602 624522
rect 306662 624456 329063 624484
rect 306662 624410 328602 624456
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 624410
rect 510007 622564 510119 622627
rect 509399 622536 510119 622564
rect 510007 621189 510119 622536
rect 510007 621077 565632 621189
rect 510005 615268 510117 615291
rect 509427 615240 510117 615268
rect 510005 614914 510117 615240
rect 510005 614802 562086 614914
rect 310208 614500 328603 614531
rect 310208 614472 329038 614500
rect 310208 614419 328603 614472
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 614419
rect 510000 607990 558540 608102
rect 510000 607972 510112 607990
rect 509383 607944 510112 607972
rect 510000 607911 510112 607944
rect 311156 604516 328600 604533
rect 311156 604488 329052 604516
rect 311156 604421 328600 604488
rect 311156 437395 311268 604421
rect 510000 600683 554994 600795
rect 510000 600676 510112 600683
rect 509371 600648 510112 600676
rect 510000 600588 510112 600648
rect 312202 594532 328600 594563
rect 312202 594504 329057 594532
rect 312202 594451 328600 594504
rect 312202 438267 312314 594451
rect 509994 593284 510106 593363
rect 509371 593256 510106 593284
rect 509994 592293 510106 593256
rect 509994 592181 551448 592293
rect 509994 585988 510106 586089
rect 509429 585960 510106 585988
rect 509994 585094 510106 585960
rect 509994 584982 547902 585094
rect 313323 584548 328616 584584
rect 313323 584520 329050 584548
rect 313323 584472 328616 584520
rect 313323 439267 313435 584472
rect 509999 578596 510111 578724
rect 509401 578568 510111 578596
rect 509999 578565 510111 578568
rect 509999 578453 544356 578565
rect 314633 574564 328599 574587
rect 314633 574536 329049 574564
rect 314633 574475 328599 574536
rect 314633 440315 314745 574475
rect 509999 571300 510111 571393
rect 509371 571283 510111 571300
rect 509371 571272 540810 571283
rect 509999 571171 540810 571272
rect 316471 564580 328600 564628
rect 316471 564552 329048 564580
rect 316471 564511 328600 564552
rect 316471 441508 316588 564511
rect 510002 564004 510114 564118
rect 509421 563976 510114 564004
rect 510002 563606 510114 563976
rect 510002 563494 537264 563606
rect 510018 556612 510130 556673
rect 509404 556584 510130 556612
rect 510018 556024 510130 556584
rect 510018 555912 533718 556024
rect 319406 554596 328603 554623
rect 319406 554568 329034 554596
rect 319406 554511 328603 554568
rect 319406 442800 319518 554511
rect 509996 549316 510108 549416
rect 509411 549288 510108 549316
rect 509996 549029 510108 549288
rect 509996 548917 530172 549029
rect 323123 544612 328604 544651
rect 323123 544584 329046 544612
rect 323123 544539 328604 544584
rect 323123 444123 323235 544539
rect 509801 542020 509913 542114
rect 509395 541992 509913 542020
rect 509801 541552 509913 541992
rect 509801 541440 526626 541552
rect 327152 534724 328633 534766
rect 509801 534724 509913 534847
rect 327152 534696 329013 534724
rect 509404 534696 509913 534724
rect 327152 534654 328633 534696
rect 327152 444904 327264 534654
rect 329005 534164 329033 534597
rect 332631 534172 332659 534627
rect 328931 534052 329388 534164
rect 332483 534060 333159 534172
rect 336257 534112 336285 534626
rect 339883 534207 339911 534610
rect 329276 445625 329388 534052
rect 333047 446277 333159 534060
rect 336122 534000 336724 534112
rect 339769 534095 340030 534207
rect 343509 534123 343537 534622
rect 347061 534198 347089 534605
rect 350687 534199 350715 534620
rect 336612 446903 336724 534000
rect 339918 447681 340030 534095
rect 343284 534011 343600 534123
rect 343284 448369 343396 534011
rect 347006 449011 347118 534198
rect 350609 534087 350815 534199
rect 354313 534100 354341 534655
rect 357939 534133 357967 534623
rect 361491 534163 361519 534624
rect 350703 449707 350815 534087
rect 353273 533988 354387 534100
rect 355959 534021 358090 534133
rect 360296 534051 361590 534163
rect 365117 534135 365145 534608
rect 368743 534142 368771 534620
rect 372369 534148 372397 534603
rect 375921 534155 375949 534636
rect 379547 534158 379575 534631
rect 353273 450523 353385 533988
rect 355959 451603 356071 534021
rect 360296 452655 360408 534051
rect 365023 534023 365488 534135
rect 368684 534030 369922 534142
rect 372278 534036 374042 534148
rect 375874 534043 378016 534155
rect 379472 534046 380597 534158
rect 383173 534135 383201 534628
rect 365376 453452 365488 534023
rect 369810 454235 369922 534030
rect 373930 454999 374042 534036
rect 377904 455774 378016 534043
rect 380485 456500 380597 534046
rect 383148 457243 383260 534135
rect 386799 534134 386827 534600
rect 385601 534022 386918 534134
rect 390351 534119 390379 534621
rect 393977 534150 394005 534608
rect 385601 458186 385713 534022
rect 388611 534007 390449 534119
rect 392644 534038 394085 534150
rect 397603 534146 397631 534646
rect 401229 534146 401257 534619
rect 388611 459251 388723 534007
rect 392644 460187 392756 534038
rect 397136 534034 397667 534146
rect 398980 534034 401393 534146
rect 404781 534138 404809 534635
rect 408407 534140 408435 534621
rect 397136 461218 397248 534034
rect 398980 462044 399092 534034
rect 403198 534026 404867 534138
rect 407350 534028 408562 534140
rect 412033 534125 412061 534617
rect 415659 534147 415687 534621
rect 419211 534174 419239 534625
rect 403198 462806 403310 534026
rect 407350 463698 407462 534028
rect 411446 534013 412164 534125
rect 415493 534035 415788 534147
rect 419127 534062 419541 534174
rect 422837 534114 422865 534607
rect 426463 534140 426491 534637
rect 430089 534151 430117 534634
rect 433715 534178 433743 534632
rect 411446 464489 411558 534013
rect 415493 465769 415605 534035
rect 419429 466884 419541 534062
rect 422788 534002 423319 534114
rect 426406 534028 427008 534140
rect 430035 534039 430556 534151
rect 433664 534066 434065 534178
rect 437267 534137 437295 534626
rect 440893 534163 440921 534638
rect 444519 534194 444547 534634
rect 423207 469267 423319 534002
rect 426896 471929 427008 534028
rect 430444 473966 430556 534039
rect 433953 476468 434065 534066
rect 437154 534025 437484 534137
rect 440817 534051 441188 534163
rect 444432 534082 444844 534194
rect 448145 534167 448173 534634
rect 437372 478866 437484 534025
rect 441076 481498 441188 534051
rect 444732 484271 444844 534082
rect 448065 534055 448497 534167
rect 451697 534145 451725 534632
rect 448385 486844 448497 534055
rect 451600 534033 451939 534145
rect 455323 534114 455351 534645
rect 458949 534148 458977 534613
rect 462575 534158 462603 534647
rect 451827 489108 451939 534033
rect 455278 534002 455600 534114
rect 458884 534036 459319 534148
rect 462500 534046 462918 534158
rect 466127 534156 466155 534624
rect 469753 534185 469781 534634
rect 455488 491118 455600 534002
rect 459207 493897 459319 534036
rect 462806 497040 462918 534046
rect 465891 534044 466231 534156
rect 469559 534072 469855 534185
rect 473379 534183 473407 534636
rect 465891 499367 466003 534044
rect 469559 501819 469672 534072
rect 473327 534071 473548 534183
rect 477005 534161 477033 534643
rect 480557 534164 480585 534628
rect 484183 534175 484211 534631
rect 473436 504226 473548 534071
rect 476959 534049 477535 534161
rect 480508 534052 481058 534164
rect 484141 534064 484976 534175
rect 487809 534156 487837 534619
rect 477423 506813 477535 534049
rect 480946 509219 481058 534052
rect 484865 511525 484976 534064
rect 487768 534044 488525 534156
rect 491435 534126 491463 534625
rect 494987 534193 495015 534621
rect 488413 513047 488525 534044
rect 491392 534014 492210 534126
rect 494929 534081 495571 534193
rect 498613 534188 498641 534626
rect 502239 534200 502267 534620
rect 505865 534200 505893 534643
rect 509417 534200 509445 534606
rect 509801 534449 509913 534696
rect 509801 534337 523080 534449
rect 492098 515275 492210 534014
rect 495459 517507 495571 534081
rect 498558 534076 500484 534188
rect 500372 520755 500484 534076
rect 502196 524032 502308 534200
rect 505820 527134 505932 534200
rect 509385 530316 509497 534200
rect 509385 530204 519534 530316
rect 505820 527022 515988 527134
rect 502196 523920 512442 524032
rect 508784 520755 508896 520811
rect 500372 520643 508896 520755
rect 495459 517395 505350 517507
rect 492098 515163 501804 515275
rect 488413 512935 498258 513047
rect 484864 511413 494712 511525
rect 480946 509107 491166 509219
rect 477423 506701 487620 506813
rect 473436 504114 484074 504226
rect 469559 501707 480528 501819
rect 465891 499255 476982 499367
rect 462806 496928 473436 497040
rect 459207 493785 469890 493897
rect 455488 491006 466344 491118
rect 451827 488996 462798 489108
rect 448385 486732 459252 486844
rect 444732 484159 455706 484271
rect 452048 481498 452160 481526
rect 441076 481386 452160 481498
rect 437372 478754 448614 478866
rect 433953 476356 445068 476468
rect 430444 473854 441522 473966
rect 426896 471817 437976 471929
rect 423207 469155 434430 469267
rect 419429 466772 430884 466884
rect 415493 465657 427338 465769
rect 411446 464377 423792 464489
rect 407350 463586 420246 463698
rect 403198 462694 416700 462806
rect 398980 461932 413154 462044
rect 409496 461218 409608 461223
rect 397136 461106 409608 461218
rect 392644 460075 406062 460187
rect 388611 459139 402516 459251
rect 385601 458074 398970 458186
rect 383148 457131 395424 457243
rect 380485 456388 391878 456500
rect 377904 455662 388332 455774
rect 373930 454887 384786 454999
rect 369810 454123 381240 454235
rect 365376 453340 377694 453452
rect 360296 452543 374148 452655
rect 355959 451491 370602 451603
rect 353273 450411 367056 450523
rect 350703 449595 363510 449707
rect 347006 448899 359964 449011
rect 343284 448257 356418 448369
rect 339918 447569 352872 447681
rect 336612 446791 349326 446903
rect 333047 446165 345780 446277
rect 329276 445513 342234 445625
rect 327152 444792 338688 444904
rect 323123 444011 335142 444123
rect 319406 442688 331596 442800
rect 316471 441396 328050 441508
rect 316471 441394 316588 441396
rect 314633 440203 324504 440315
rect 313323 439155 320958 439267
rect 312202 438155 317412 438267
rect 311156 437283 313866 437395
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 437283
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 438155
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 439155
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 440203
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 441396
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 442688
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 444011
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 444792
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 445513
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 446165
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 446791
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 447569
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 448257
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 448899
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 449595
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 450411
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 451491
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 452543
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 453340
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 454123
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 454887
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 455662
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 456388
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 457131
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 458074
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 459139
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 460075
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 461106
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 461932
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 462694
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 463586
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 464377
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 465657
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 466772
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 469155
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 471817
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 473854
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 476356
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 478754
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 481386
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 484159
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 486732
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 488996
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 491006
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 493785
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 496928
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 499255
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 501707
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 504114
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 506701
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 509107
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 511413
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 512935
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 515163
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 517395
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 520643
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 523920
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 527022
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 530204
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 534337
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 541440
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 548917
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 555912
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 563494
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 571171
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 578453
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 584982
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 592181
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 600683
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 607990
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 614802
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 621077
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 629319
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 637291
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 644144
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 120805 690305 124595 694095
rect 68805 673405 72395 676995
rect 16812 658612 20388 662188
rect 414005 693505 417795 697295
rect 466005 696905 469795 700695
rect 567208 687508 570992 691292
rect 573705 678405 577895 682595
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 16800 700000 20400 702300
rect -800 680242 1700 685242
rect 16807 662188 20393 700000
rect 68800 676995 72400 702300
rect 120800 694095 124600 702300
rect 120800 690305 120805 694095
rect 124595 690305 124600 694095
rect 414000 697295 417800 702300
rect 414000 693505 414005 697295
rect 417795 693505 417800 697295
rect 466000 700695 469800 702300
rect 466000 696905 466005 700695
rect 469795 696905 469800 700695
rect 567200 700600 571000 702300
rect 466000 696900 469800 696905
rect 414000 693500 417800 693505
rect 120800 690300 124600 690305
rect 567203 691292 570997 700600
rect 567203 687508 567208 691292
rect 570992 687508 570997 691292
rect 567203 687503 570997 687508
rect 582300 682600 584800 682984
rect 573700 682595 584800 682600
rect 573700 678405 573705 682595
rect 577895 678405 584800 682595
rect 573700 678400 584800 678405
rect 582300 677984 584800 678400
rect 68800 673405 68805 676995
rect 72395 673405 72400 676995
rect 68800 673400 72400 673405
rect 16807 658612 16812 662188
rect 20388 658612 20393 662188
rect 16807 658607 20393 658612
rect -800 643842 298770 648642
rect 301230 643842 301236 648642
rect 307588 643566 313656 650884
rect 527956 643566 534024 650946
rect 307588 643366 329182 643566
rect 509268 643366 534024 643566
rect 307588 641166 313656 643366
rect 327770 642366 327970 642372
rect 327970 642166 329182 642366
rect 509268 642166 510096 642366
rect 510296 642166 510302 642366
rect 327770 642160 327970 642166
rect 527956 641166 534024 643366
rect 578106 642244 578436 644584
rect 307588 640966 329182 641166
rect 509268 640966 534024 641166
rect 307588 638766 313656 640966
rect 327764 639766 327770 639966
rect 327970 639766 329182 639966
rect 509268 639766 510092 639966
rect 510292 639766 510298 639966
rect 527956 638766 534024 640966
rect 569598 639784 569604 642244
rect 572064 642124 578436 642244
rect 580896 642124 584800 644584
rect 572064 639784 584800 642124
rect -800 633842 298770 638642
rect 301230 633842 301236 638642
rect 307588 638566 329182 638766
rect 509268 638566 534024 638766
rect 307588 636366 313656 638566
rect 327762 637366 327768 637566
rect 327968 637366 329182 637566
rect 509268 637366 510084 637566
rect 510284 637366 510290 637566
rect 527956 636366 534024 638566
rect 307588 636166 329182 636366
rect 509268 636166 534024 636366
rect 307588 633966 313656 636166
rect 327782 634966 327788 635166
rect 327988 634966 329182 635166
rect 509268 634966 510100 635166
rect 510300 634966 510306 635166
rect 527956 633966 534024 636166
rect 307588 633766 329182 633966
rect 509268 633766 534024 633966
rect 307588 631566 313656 633766
rect 327794 632566 327800 632766
rect 328000 632566 329182 632766
rect 509268 632566 510108 632766
rect 510308 632566 510314 632766
rect 527956 631566 534024 633766
rect 572598 632124 572604 634584
rect 575064 632244 584800 634584
rect 575064 632124 576894 632244
rect 307588 631366 329182 631566
rect 509268 631366 534024 631566
rect 307588 629166 313656 631366
rect 327774 630166 327780 630366
rect 327980 630166 329182 630366
rect 509268 630166 510114 630366
rect 510314 630166 510320 630366
rect 527956 629166 534024 631366
rect 576888 629784 576894 632124
rect 579354 629784 584800 632244
rect 307588 628966 329182 629166
rect 509268 628966 534024 629166
rect 307588 626766 313656 628966
rect 327758 627766 327764 627966
rect 327964 627766 329182 627966
rect 509268 627766 510106 627966
rect 510306 627766 510312 627966
rect 527956 626766 534024 628966
rect 307588 626566 329182 626766
rect 509268 626566 534024 626766
rect 307588 624366 313656 626566
rect 327772 625366 327778 625566
rect 327978 625366 329182 625566
rect 509268 625366 510114 625566
rect 510314 625366 510320 625566
rect 527956 624366 534024 626566
rect 307588 624166 329182 624366
rect 509268 624166 534024 624366
rect 307588 621966 313656 624166
rect 327772 622966 327778 623166
rect 327978 622966 329182 623166
rect 509268 622966 510112 623166
rect 510312 622966 510318 623166
rect 527956 621966 534024 624166
rect 307588 621766 329182 621966
rect 509268 621766 534024 621966
rect 307588 619566 313656 621766
rect 327780 620566 327786 620766
rect 327986 620566 329182 620766
rect 509268 620566 510114 620766
rect 510314 620566 510320 620766
rect 527956 619566 534024 621766
rect 307588 619366 329182 619566
rect 509268 619366 534024 619566
rect 307588 617166 313656 619366
rect 327786 618166 327792 618366
rect 327992 618166 329182 618366
rect 509268 618166 510106 618366
rect 510306 618166 510312 618366
rect 527956 617166 534024 619366
rect 307588 616966 329182 617166
rect 509268 616966 534024 617166
rect 307588 614766 313656 616966
rect 327804 615766 327810 615966
rect 328010 615766 329182 615966
rect 509268 615766 510106 615966
rect 510306 615766 510312 615966
rect 307588 614566 329182 614766
rect 307588 610382 313656 614566
rect 327816 613366 327822 613566
rect 328022 613366 329182 613566
rect 509268 613366 510128 613566
rect 510328 613366 510334 613566
rect 327822 611382 327828 611582
rect 328028 611382 329182 611582
rect 509268 611382 510136 611582
rect 510336 611382 510342 611582
rect 527956 610382 534024 616966
rect 307588 610182 329182 610382
rect 509268 610182 534024 610382
rect 307588 607982 313656 610182
rect 327838 608982 327844 609182
rect 328044 608982 329182 609182
rect 509268 608982 510146 609182
rect 510346 608982 510352 609182
rect 527956 607982 534024 610182
rect 307588 607782 329182 607982
rect 509268 607782 534024 607982
rect 307588 605582 313656 607782
rect 327844 606582 327850 606782
rect 328050 606582 329182 606782
rect 509268 606582 510150 606782
rect 510350 606582 510356 606782
rect 527956 605582 534024 607782
rect 307588 605382 329182 605582
rect 509268 605382 534024 605582
rect 307588 603182 313656 605382
rect 327852 604182 327858 604382
rect 328058 604182 329182 604382
rect 509268 604182 510136 604382
rect 510336 604182 510342 604382
rect 527956 603182 534024 605382
rect 307588 602982 329182 603182
rect 509268 602982 534024 603182
rect 307588 600782 313656 602982
rect 327858 601782 327864 601982
rect 328064 601782 329182 601982
rect 509268 601782 510138 601982
rect 510338 601782 510344 601982
rect 527956 600782 534024 602982
rect 307588 600582 329182 600782
rect 509268 600582 534024 600782
rect 307588 598724 313656 600582
rect 327884 599382 327890 599582
rect 328090 599382 329182 599582
rect 509268 599382 510130 599582
rect 510330 599382 510336 599582
rect 327600 598724 327800 598800
rect 307588 598723 327800 598724
rect 307588 598325 327341 598723
rect 327739 598600 327800 598723
rect 516317 598600 516715 598605
rect 527956 598600 534024 600582
rect 327739 598500 327740 598600
rect 516316 598599 534024 598600
rect 327739 598325 327800 598500
rect 307588 598324 327800 598325
rect 307588 595414 313656 598324
rect 327600 598300 327800 598324
rect 516316 598201 516317 598599
rect 516715 598201 534024 598599
rect 516316 598200 534024 598201
rect 516317 598195 516715 598200
rect 327870 596214 327876 596414
rect 328076 596214 329182 596414
rect 328100 595414 328300 595500
rect 307588 595413 328300 595414
rect 307588 595015 327813 595413
rect 328211 595300 328300 595413
rect 510300 595414 510500 595500
rect 527956 595414 534024 598200
rect 510300 595413 534024 595414
rect 510300 595300 510461 595413
rect 328211 595200 328212 595300
rect 328211 595015 328300 595200
rect 510460 595100 510461 595300
rect 307588 595014 328300 595015
rect 307588 593198 313656 595014
rect 328100 595000 328300 595014
rect 510300 595015 510461 595100
rect 510859 595015 534024 595413
rect 510300 595014 534024 595015
rect 510300 594900 510500 595014
rect 327912 594198 327918 594398
rect 328118 594198 329182 594398
rect 509268 594198 510568 594398
rect 510768 594198 510774 594398
rect 527956 593198 534024 595014
rect 307588 592998 329182 593198
rect 509268 592998 534024 593198
rect 307588 591414 313656 592998
rect 327934 591798 327940 591998
rect 328140 591798 329182 591998
rect 509268 591798 510568 591998
rect 510768 591798 510774 591998
rect 327900 591414 328100 591500
rect 307588 591413 328100 591414
rect 307588 591015 327693 591413
rect 328091 591300 328100 591413
rect 510300 591414 510500 591500
rect 527956 591414 534024 592998
rect 510300 591413 534024 591414
rect 510300 591300 510423 591413
rect 328091 591200 328092 591300
rect 328091 591015 328100 591200
rect 510422 591100 510423 591300
rect 307588 591014 328100 591015
rect 307588 590798 313656 591014
rect 327900 591000 328100 591014
rect 510300 591015 510423 591100
rect 510821 591015 534024 591413
rect 510300 591014 534024 591015
rect 510300 590900 510500 591014
rect 527956 590798 534024 591014
rect 307588 590598 329182 590798
rect 509268 590598 534024 590798
rect 307588 588398 313656 590598
rect 327948 589398 327954 589598
rect 328154 589398 329182 589598
rect 509268 589398 510560 589598
rect 510760 589398 510766 589598
rect 527956 588398 534024 590598
rect 583520 589472 584800 589584
rect 307588 588198 329182 588398
rect 509268 588198 534024 588398
rect 583520 588290 584800 588402
rect 307588 587414 313656 588198
rect 327600 587414 327800 587500
rect 307588 587413 327800 587414
rect 307588 587015 327345 587413
rect 327743 587300 327800 587413
rect 511000 587414 511200 587500
rect 527956 587414 534024 588198
rect 511000 587413 534024 587414
rect 511000 587300 511099 587413
rect 327743 587200 327744 587300
rect 327743 587015 327800 587200
rect 307588 587014 327800 587015
rect 307588 585998 313656 587014
rect 327600 587000 327800 587014
rect 328020 586998 329182 587198
rect 509268 586998 510462 587198
rect 511098 587100 511099 587300
rect 328020 586614 328220 586998
rect 510262 586818 510462 586998
rect 511000 587015 511099 587100
rect 511497 587015 534024 587413
rect 583520 587108 584800 587220
rect 511000 587014 534024 587015
rect 511000 586900 511200 587014
rect 510256 586618 510262 586818
rect 510462 586618 510468 586818
rect 326864 586414 326870 586614
rect 327070 586414 328220 586614
rect 527956 585998 534024 587014
rect 307588 585798 329182 585998
rect 509268 585798 534024 585998
rect 583520 585926 584800 586038
rect 307588 583598 313656 585798
rect 326868 584598 326874 584798
rect 327074 584598 329182 584798
rect 509268 584598 510280 584798
rect 510480 584598 510486 584798
rect 527956 583598 534024 585798
rect 583520 584744 584800 584856
rect 307588 583413 329182 583598
rect 307588 583015 327855 583413
rect 328253 583398 329182 583413
rect 509268 583413 534024 583598
rect 583520 583562 584800 583674
rect 509268 583398 510449 583413
rect 328253 583200 328254 583398
rect 328253 583015 328400 583200
rect 510448 583100 510449 583398
rect 307588 583014 328400 583015
rect 307588 580814 313656 583014
rect 328200 583000 328400 583014
rect 510300 583015 510449 583100
rect 510847 583015 534024 583413
rect 510300 583014 534024 583015
rect 510300 582900 510500 583014
rect 326878 582198 326884 582398
rect 327084 582198 329182 582398
rect 509268 582198 510548 582398
rect 510748 582198 510754 582398
rect 307588 580614 329182 580814
rect 307588 578714 313656 580614
rect 326866 579414 326872 579614
rect 327072 579414 329182 579614
rect 510300 579414 510500 579500
rect 527956 579414 534024 583014
rect 510300 579413 534024 579414
rect 510300 579300 510441 579413
rect 510440 579100 510441 579300
rect 510300 579015 510441 579100
rect 510839 579015 534024 579413
rect 510300 579014 534024 579015
rect 510300 578900 510500 579014
rect 327483 578714 327881 578719
rect 307588 578713 327882 578714
rect 307588 578315 327483 578713
rect 327881 578400 327882 578713
rect 327881 578315 328000 578400
rect 307588 578314 328000 578315
rect 307588 576014 313656 578314
rect 327483 578309 328000 578314
rect 327800 578200 328000 578309
rect 326884 577014 326890 577214
rect 327090 577014 329182 577214
rect 509268 577014 510542 577214
rect 510742 577014 510748 577214
rect 527956 576014 534024 579014
rect 307588 575814 329182 576014
rect 509268 575814 534024 576014
rect 307588 575414 313656 575814
rect 327800 575414 328000 575500
rect 307588 575413 328000 575414
rect 307588 575015 327441 575413
rect 327839 575300 328000 575413
rect 510400 575414 510600 575500
rect 527956 575414 534024 575814
rect 510400 575413 534024 575414
rect 510400 575300 510487 575413
rect 327839 575200 327840 575300
rect 327839 575015 328000 575200
rect 510486 575100 510487 575300
rect 307588 575014 328000 575015
rect 307588 573614 313656 575014
rect 327800 575000 328000 575014
rect 510400 575015 510487 575100
rect 510885 575015 534024 575413
rect 510400 575014 534024 575015
rect 510400 574900 510600 575014
rect 327568 574614 327574 574814
rect 327774 574614 329182 574814
rect 509268 574614 510548 574814
rect 510748 574614 510754 574814
rect 527956 573614 534024 575014
rect 307588 573414 329182 573614
rect 509268 573414 534024 573614
rect 307588 571414 313656 573414
rect 327570 572214 327576 572414
rect 327776 572214 329182 572414
rect 509268 572214 510542 572414
rect 510742 572214 510748 572414
rect 327800 571414 328000 571500
rect 307588 571413 328000 571414
rect 307588 571015 327511 571413
rect 327909 571300 328000 571413
rect 510300 571414 510600 571500
rect 527956 571414 534024 573414
rect 510300 571413 534024 571414
rect 510300 571300 510433 571413
rect 327909 571214 327910 571300
rect 510432 571214 510433 571300
rect 327909 571015 329182 571214
rect 307588 571014 329182 571015
rect 509268 571015 510433 571214
rect 510831 571015 534024 571413
rect 509268 571014 534024 571015
rect 307588 568814 313656 571014
rect 327604 569814 327610 570014
rect 327810 569814 329182 570014
rect 509268 569814 510520 570014
rect 510720 569814 510726 570014
rect 527956 568814 534024 571014
rect 307588 568614 329182 568814
rect 509268 568614 534024 568814
rect 307588 567152 313656 568614
rect 327620 567414 327626 567614
rect 327826 567414 329182 567614
rect 509268 567414 510520 567614
rect 510720 567414 510726 567614
rect 326837 567152 327235 567157
rect 307588 567151 327236 567152
rect 307588 566753 326837 567151
rect 327235 566753 327236 567151
rect 510800 567130 511000 567200
rect 527956 567130 534024 568614
rect 510800 567129 534024 567130
rect 510800 567000 510895 567129
rect 510894 566800 510895 567000
rect 307588 566752 327236 566753
rect 307588 566414 313656 566752
rect 326837 566747 327235 566752
rect 510800 566731 510895 566800
rect 511293 566731 534024 567129
rect 510800 566730 534024 566731
rect 510800 566600 511000 566730
rect 527956 566414 534024 566730
rect 307588 566214 329182 566414
rect 509268 566214 534024 566414
rect -800 559442 1660 564242
rect 307588 558830 313656 566214
rect 327610 565014 327616 565214
rect 327816 565014 329182 565214
rect 509268 565014 510542 565214
rect 510742 565014 510748 565214
rect 510632 560030 510832 560036
rect 327234 559830 327240 560030
rect 327440 559830 329182 560030
rect 509268 559830 510632 560030
rect 510632 559824 510832 559830
rect 527956 558830 534024 566214
rect 307588 558630 329182 558830
rect 509268 558630 534024 558830
rect 307588 556430 313656 558630
rect 327234 557630 327434 557636
rect 327434 557430 329182 557630
rect 509268 557430 510646 557630
rect 510846 557430 510852 557630
rect 327234 557424 327434 557430
rect 527956 556430 534024 558630
rect 307588 556230 329182 556430
rect 509268 556230 534024 556430
rect -800 549442 1660 554242
rect 307588 554030 313656 556230
rect 327228 555030 327234 555230
rect 327434 555030 329182 555230
rect 509268 555030 510628 555230
rect 510828 555030 510834 555230
rect 527956 554030 534024 556230
rect 307588 553830 329182 554030
rect 509268 553830 534024 554030
rect 307588 551630 313656 553830
rect 327232 552630 327238 552830
rect 327438 552630 329182 552830
rect 509268 552630 510624 552830
rect 510824 552630 510830 552830
rect 527956 551630 534024 553830
rect 307588 551430 329182 551630
rect 509268 551430 534024 551630
rect 307588 549230 313656 551430
rect 327212 550230 327218 550430
rect 327418 550230 329182 550430
rect 509268 550230 510618 550430
rect 510818 550230 510824 550430
rect 527956 549230 534024 551430
rect 582340 550562 584800 555362
rect 307588 549030 329182 549230
rect 509268 549030 534024 549230
rect 307588 526210 313656 549030
rect 510606 548030 510806 548036
rect 327214 547830 327220 548030
rect 327420 547830 329182 548030
rect 509268 547830 510606 548030
rect 510606 547824 510806 547830
rect 527956 526210 534024 549030
rect 582340 540562 584800 545362
rect 307442 520142 534024 526210
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 307588 196230 313656 520142
rect 331170 196230 335970 520142
rect 352630 196230 357430 520142
rect 375779 196230 380582 520142
rect 403950 196230 408750 520142
rect 428378 196230 433182 520142
rect 457269 196230 462071 520142
rect 484680 196230 489480 520142
rect 523110 196230 527910 520142
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 288040 191430 584800 196230
rect 331170 186230 335970 191430
rect 375779 186230 380582 191430
rect 428378 186230 433182 191430
rect 457269 191429 462071 191430
rect 484680 186230 489480 191430
rect 288040 181430 584800 186230
rect 375779 181429 380582 181430
rect 428378 181428 433182 181430
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 298770 643842 301230 648642
rect 327770 642166 327970 642366
rect 510096 642166 510296 642366
rect 327770 639766 327970 639966
rect 510092 639766 510292 639966
rect 569604 639784 572064 642244
rect 578436 642124 580896 644584
rect 298770 633842 301230 638642
rect 327768 637366 327968 637566
rect 510084 637366 510284 637566
rect 327788 634966 327988 635166
rect 510100 634966 510300 635166
rect 327800 632566 328000 632766
rect 510108 632566 510308 632766
rect 572604 632124 575064 634584
rect 327780 630166 327980 630366
rect 510114 630166 510314 630366
rect 576894 629784 579354 632244
rect 327764 627766 327964 627966
rect 510106 627766 510306 627966
rect 327778 625366 327978 625566
rect 510114 625366 510314 625566
rect 327778 622966 327978 623166
rect 510112 622966 510312 623166
rect 327786 620566 327986 620766
rect 510114 620566 510314 620766
rect 327792 618166 327992 618366
rect 510106 618166 510306 618366
rect 327810 615766 328010 615966
rect 510106 615766 510306 615966
rect 327822 613366 328022 613566
rect 510128 613366 510328 613566
rect 327828 611382 328028 611582
rect 510136 611382 510336 611582
rect 327844 608982 328044 609182
rect 510146 608982 510346 609182
rect 327850 606582 328050 606782
rect 510150 606582 510350 606782
rect 327858 604182 328058 604382
rect 510136 604182 510336 604382
rect 327864 601782 328064 601982
rect 510138 601782 510338 601982
rect 327890 599382 328090 599582
rect 510130 599382 510330 599582
rect 327341 598325 327739 598723
rect 516317 598201 516715 598599
rect 327876 596214 328076 596414
rect 327813 595015 328211 595413
rect 510461 595015 510859 595413
rect 327918 594198 328118 594398
rect 510568 594198 510768 594398
rect 327940 591798 328140 591998
rect 510568 591798 510768 591998
rect 327693 591015 328091 591413
rect 510423 591015 510821 591413
rect 327954 589398 328154 589598
rect 510560 589398 510760 589598
rect 327345 587015 327743 587413
rect 511099 587015 511497 587413
rect 510262 586618 510462 586818
rect 326870 586414 327070 586614
rect 326874 584598 327074 584798
rect 510280 584598 510480 584798
rect 327855 583015 328253 583413
rect 510449 583015 510847 583413
rect 326884 582198 327084 582398
rect 510548 582198 510748 582398
rect 326872 579414 327072 579614
rect 510441 579015 510839 579413
rect 327483 578315 327881 578713
rect 326890 577014 327090 577214
rect 510542 577014 510742 577214
rect 327441 575015 327839 575413
rect 510487 575015 510885 575413
rect 327574 574614 327774 574814
rect 510548 574614 510748 574814
rect 327576 572214 327776 572414
rect 510542 572214 510742 572414
rect 327511 571015 327909 571413
rect 510433 571015 510831 571413
rect 327610 569814 327810 570014
rect 510520 569814 510720 570014
rect 327626 567414 327826 567614
rect 510520 567414 510720 567614
rect 326837 566753 327235 567151
rect 510895 566731 511293 567129
rect 327616 565014 327816 565214
rect 510542 565014 510742 565214
rect 327240 559830 327440 560030
rect 510632 559830 510832 560030
rect 327234 557430 327434 557630
rect 510646 557430 510846 557630
rect 327234 555030 327434 555230
rect 510628 555030 510828 555230
rect 327238 552630 327438 552830
rect 510624 552630 510824 552830
rect 327218 550230 327418 550430
rect 510618 550230 510818 550430
rect 327220 547830 327420 548030
rect 510606 547830 510806 548030
<< metal4 >>
rect 297340 648642 303408 650884
rect 297340 643842 298770 648642
rect 301230 643842 303408 648642
rect 297340 642366 303408 643842
rect 327769 642366 327971 642367
rect 297340 642166 327770 642366
rect 327970 642166 327971 642366
rect 297340 639966 303408 642166
rect 327769 642165 327971 642166
rect 510095 642366 510297 642367
rect 537254 642366 543322 650924
rect 510095 642166 510096 642366
rect 510296 642166 543322 642366
rect 580895 644584 580897 644585
rect 510095 642165 510297 642166
rect 327769 639966 327971 639967
rect 297340 639766 327770 639966
rect 327970 639766 327971 639966
rect 297340 638642 303408 639766
rect 327769 639765 327971 639766
rect 510091 639966 510293 639967
rect 537254 639966 543322 642166
rect 510091 639766 510092 639966
rect 510292 639766 543322 639966
rect 580896 642124 580897 644584
rect 580895 642123 580897 642124
rect 510091 639765 510293 639766
rect 297340 633842 298770 638642
rect 301230 637566 303408 638642
rect 327767 637566 327969 637567
rect 301230 637366 327768 637566
rect 327968 637366 327969 637566
rect 301230 635166 303408 637366
rect 327767 637365 327969 637366
rect 510083 637566 510285 637567
rect 537254 637566 543322 639766
rect 510083 637366 510084 637566
rect 510284 637366 543322 637566
rect 510083 637365 510285 637366
rect 327787 635166 327989 635167
rect 301230 634966 327788 635166
rect 327988 634966 327989 635166
rect 301230 633842 303408 634966
rect 327787 634965 327989 634966
rect 510099 635166 510301 635167
rect 537254 635166 543322 637366
rect 510099 634966 510100 635166
rect 510300 634966 543322 635166
rect 510099 634965 510301 634966
rect 297340 632766 303408 633842
rect 327799 632766 328001 632767
rect 297340 632566 327800 632766
rect 328000 632566 328001 632766
rect 297340 630366 303408 632566
rect 327799 632565 328001 632566
rect 510107 632766 510309 632767
rect 537254 632766 543322 634966
rect 510107 632566 510108 632766
rect 510308 632566 543322 632766
rect 510107 632565 510309 632566
rect 327779 630366 327981 630367
rect 297340 630166 327780 630366
rect 327980 630166 327981 630366
rect 297340 627966 303408 630166
rect 327779 630165 327981 630166
rect 510113 630366 510315 630367
rect 537254 630366 543322 632566
rect 575063 634584 575065 634585
rect 575064 632124 575065 634584
rect 575063 632123 575065 632124
rect 579353 632244 579355 632245
rect 510113 630166 510114 630366
rect 510314 630166 543322 630366
rect 510113 630165 510315 630166
rect 327763 627966 327965 627967
rect 297340 627766 327764 627966
rect 327964 627766 327965 627966
rect 297340 625566 303408 627766
rect 327763 627765 327965 627766
rect 510105 627966 510307 627967
rect 537254 627966 543322 630166
rect 579354 629784 579355 632244
rect 579353 629783 579355 629784
rect 510105 627766 510106 627966
rect 510306 627766 543322 627966
rect 510105 627765 510307 627766
rect 327777 625566 327979 625567
rect 297340 625366 327778 625566
rect 327978 625366 327979 625566
rect 297340 623166 303408 625366
rect 327777 625365 327979 625366
rect 510113 625566 510315 625567
rect 537254 625566 543322 627766
rect 510113 625366 510114 625566
rect 510314 625366 543322 625566
rect 510113 625365 510315 625366
rect 327777 623166 327979 623167
rect 297340 622966 327778 623166
rect 327978 622966 327979 623166
rect 297340 620766 303408 622966
rect 327777 622965 327979 622966
rect 510111 623166 510313 623167
rect 537254 623166 543322 625366
rect 510111 622966 510112 623166
rect 510312 622966 543322 623166
rect 510111 622965 510313 622966
rect 327785 620766 327987 620767
rect 297340 620566 327786 620766
rect 327986 620566 327987 620766
rect 297340 618366 303408 620566
rect 327785 620565 327987 620566
rect 510113 620766 510315 620767
rect 537254 620766 543322 622966
rect 510113 620566 510114 620766
rect 510314 620566 543322 620766
rect 510113 620565 510315 620566
rect 327791 618366 327993 618367
rect 297340 618166 327792 618366
rect 327992 618166 327993 618366
rect 297340 615966 303408 618166
rect 327791 618165 327993 618166
rect 510105 618366 510307 618367
rect 537254 618366 543322 620566
rect 510105 618166 510106 618366
rect 510306 618166 543322 618366
rect 510105 618165 510307 618166
rect 327809 615966 328011 615967
rect 297340 615766 327810 615966
rect 328010 615766 328011 615966
rect 297340 613566 303408 615766
rect 327809 615765 328011 615766
rect 510105 615966 510307 615967
rect 537254 615966 543322 618166
rect 510105 615766 510106 615966
rect 510306 615766 543322 615966
rect 510105 615765 510307 615766
rect 327821 613566 328023 613567
rect 297340 613366 327822 613566
rect 328022 613366 328023 613566
rect 297340 611582 303408 613366
rect 327821 613365 328023 613366
rect 510127 613566 510329 613567
rect 537254 613566 543322 615766
rect 510127 613366 510128 613566
rect 510328 613366 543322 613566
rect 510127 613365 510329 613366
rect 327827 611582 328029 611583
rect 297340 611382 327828 611582
rect 328028 611382 328029 611582
rect 297340 609182 303408 611382
rect 327827 611381 328029 611382
rect 510135 611582 510337 611583
rect 537254 611582 543322 613366
rect 510135 611382 510136 611582
rect 510336 611382 543322 611582
rect 510135 611381 510337 611382
rect 327843 609182 328045 609183
rect 297340 608982 327844 609182
rect 328044 608982 328045 609182
rect 297340 606782 303408 608982
rect 327843 608981 328045 608982
rect 510145 609182 510347 609183
rect 537254 609182 543322 611382
rect 510145 608982 510146 609182
rect 510346 608982 543322 609182
rect 510145 608981 510347 608982
rect 327849 606782 328051 606783
rect 297340 606582 327850 606782
rect 328050 606582 328051 606782
rect 297340 604382 303408 606582
rect 327849 606581 328051 606582
rect 510149 606782 510351 606783
rect 537254 606782 543322 608982
rect 510149 606582 510150 606782
rect 510350 606582 543322 606782
rect 510149 606581 510351 606582
rect 327857 604382 328059 604383
rect 297340 604182 327858 604382
rect 328058 604182 328059 604382
rect 297340 601982 303408 604182
rect 327857 604181 328059 604182
rect 510135 604382 510337 604383
rect 537254 604382 543322 606582
rect 510135 604182 510136 604382
rect 510336 604182 543322 604382
rect 510135 604181 510337 604182
rect 327863 601982 328065 601983
rect 297340 601782 327864 601982
rect 328064 601782 328065 601982
rect 297340 599582 303408 601782
rect 327863 601781 328065 601782
rect 510137 601982 510339 601983
rect 537254 601982 543322 604182
rect 510137 601782 510138 601982
rect 510338 601782 543322 601982
rect 510137 601781 510339 601782
rect 327889 599582 328091 599583
rect 297340 599382 327890 599582
rect 328090 599382 328091 599582
rect 297340 596414 303408 599382
rect 327889 599381 328091 599382
rect 510129 599582 510331 599583
rect 537254 599582 543322 601782
rect 510129 599382 510130 599582
rect 510330 599382 543322 599582
rect 510129 599381 510331 599382
rect 327340 598723 327740 598724
rect 327340 598325 327341 598723
rect 327739 598325 327740 598723
rect 327340 598324 327740 598325
rect 516316 598599 516716 598600
rect 516316 598201 516317 598599
rect 516715 598201 516716 598599
rect 516316 598200 516716 598201
rect 327875 596414 328077 596415
rect 297340 596214 327876 596414
rect 328076 596214 328077 596414
rect 297340 594398 303408 596214
rect 327875 596213 328077 596214
rect 327812 595413 328212 595414
rect 327812 595015 327813 595413
rect 328211 595015 328212 595413
rect 327812 595014 328212 595015
rect 510460 595413 510860 595414
rect 510460 595015 510461 595413
rect 510859 595015 510860 595413
rect 510460 595014 510860 595015
rect 327917 594398 328119 594399
rect 297340 594198 327918 594398
rect 328118 594198 328119 594398
rect 297340 591998 303408 594198
rect 327917 594197 328119 594198
rect 510567 594398 510769 594399
rect 537254 594398 543322 599382
rect 510567 594198 510568 594398
rect 510768 594198 543322 594398
rect 510567 594197 510769 594198
rect 327939 591998 328141 591999
rect 297340 591798 327940 591998
rect 328140 591798 328141 591998
rect 297340 589598 303408 591798
rect 327939 591797 328141 591798
rect 510567 591998 510769 591999
rect 537254 591998 543322 594198
rect 510567 591798 510568 591998
rect 510768 591798 543322 591998
rect 510567 591797 510769 591798
rect 327692 591413 328092 591414
rect 327692 591015 327693 591413
rect 328091 591015 328092 591413
rect 327692 591014 328092 591015
rect 510422 591413 510822 591414
rect 510422 591015 510423 591413
rect 510821 591015 510822 591413
rect 510422 591014 510822 591015
rect 327953 589598 328155 589599
rect 297340 589398 327954 589598
rect 328154 589398 328155 589598
rect 297340 586614 303408 589398
rect 327953 589397 328155 589398
rect 510559 589598 510761 589599
rect 537254 589598 543322 591798
rect 510559 589398 510560 589598
rect 510760 589398 543322 589598
rect 510559 589397 510761 589398
rect 327344 587413 327744 587414
rect 327344 587015 327345 587413
rect 327743 587015 327744 587413
rect 327344 587014 327744 587015
rect 511098 587413 511498 587414
rect 511098 587015 511099 587413
rect 511497 587015 511498 587413
rect 511098 587014 511498 587015
rect 510261 586818 510463 586819
rect 537254 586818 543322 589398
rect 510261 586618 510262 586818
rect 510462 586618 543322 586818
rect 510261 586617 510463 586618
rect 326869 586614 327071 586615
rect 297340 586414 326870 586614
rect 327070 586414 327071 586614
rect 297340 584798 303408 586414
rect 326869 586413 327071 586414
rect 326873 584798 327075 584799
rect 297340 584598 326874 584798
rect 327074 584598 327075 584798
rect 297340 582398 303408 584598
rect 326873 584597 327075 584598
rect 510279 584798 510481 584799
rect 537254 584798 543322 586618
rect 510279 584598 510280 584798
rect 510480 584598 543322 584798
rect 510279 584597 510481 584598
rect 327854 583413 328254 583414
rect 327854 583015 327855 583413
rect 328253 583015 328254 583413
rect 327854 583014 328254 583015
rect 510448 583413 510848 583414
rect 510448 583015 510449 583413
rect 510847 583015 510848 583413
rect 510448 583014 510848 583015
rect 326883 582398 327085 582399
rect 297340 582198 326884 582398
rect 327084 582198 327085 582398
rect 297340 579614 303408 582198
rect 326883 582197 327085 582198
rect 510547 582398 510749 582399
rect 537254 582398 543322 584598
rect 510547 582198 510548 582398
rect 510748 582198 543322 582398
rect 510547 582197 510749 582198
rect 326871 579614 327073 579615
rect 297340 579414 326872 579614
rect 327072 579414 327073 579614
rect 297340 577214 303408 579414
rect 326871 579413 327073 579414
rect 510440 579413 510840 579414
rect 510440 579015 510441 579413
rect 510839 579015 510840 579413
rect 510440 579014 510840 579015
rect 327482 578713 327882 578714
rect 327482 578315 327483 578713
rect 327881 578315 327882 578713
rect 327482 578314 327882 578315
rect 326889 577214 327091 577215
rect 297340 577014 326890 577214
rect 327090 577014 327091 577214
rect 297340 574814 303408 577014
rect 326889 577013 327091 577014
rect 510541 577214 510743 577215
rect 537254 577214 543322 582198
rect 510541 577014 510542 577214
rect 510742 577014 543322 577214
rect 510541 577013 510743 577014
rect 327440 575413 327840 575414
rect 327440 575015 327441 575413
rect 327839 575015 327840 575413
rect 327440 575014 327840 575015
rect 510486 575413 510886 575414
rect 510486 575015 510487 575413
rect 510885 575015 510886 575413
rect 510486 575014 510886 575015
rect 327573 574814 327775 574815
rect 297340 574614 327574 574814
rect 327774 574614 327775 574814
rect 297340 572414 303408 574614
rect 327573 574613 327775 574614
rect 510547 574814 510749 574815
rect 537254 574814 543322 577014
rect 510547 574614 510548 574814
rect 510748 574614 543322 574814
rect 510547 574613 510749 574614
rect 327575 572414 327777 572415
rect 297340 572214 327576 572414
rect 327776 572214 327777 572414
rect 297340 570014 303408 572214
rect 327575 572213 327777 572214
rect 510541 572414 510743 572415
rect 537254 572414 543322 574614
rect 510541 572214 510542 572414
rect 510742 572214 543322 572414
rect 510541 572213 510743 572214
rect 327510 571413 327910 571414
rect 327510 571015 327511 571413
rect 327909 571015 327910 571413
rect 327510 571014 327910 571015
rect 510432 571413 510832 571414
rect 510432 571015 510433 571413
rect 510831 571015 510832 571413
rect 510432 571014 510832 571015
rect 327609 570014 327811 570015
rect 297340 569814 327610 570014
rect 327810 569814 327811 570014
rect 297340 567614 303408 569814
rect 327609 569813 327811 569814
rect 510519 570014 510721 570015
rect 537254 570014 543322 572214
rect 510519 569814 510520 570014
rect 510720 569814 543322 570014
rect 510519 569813 510721 569814
rect 327625 567614 327827 567615
rect 297340 567414 327626 567614
rect 327826 567414 327827 567614
rect 297340 565214 303408 567414
rect 327625 567413 327827 567414
rect 510519 567614 510721 567615
rect 537254 567614 543322 569814
rect 510519 567414 510520 567614
rect 510720 567414 543322 567614
rect 510519 567413 510721 567414
rect 326836 567151 327236 567152
rect 326836 566753 326837 567151
rect 327235 566753 327236 567151
rect 326836 566752 327236 566753
rect 510894 567129 511294 567130
rect 510894 566731 510895 567129
rect 511293 566731 511294 567129
rect 510894 566730 511294 566731
rect 327615 565214 327817 565215
rect 297340 565014 327616 565214
rect 327816 565014 327817 565214
rect 297340 560030 303408 565014
rect 327615 565013 327817 565014
rect 510541 565214 510743 565215
rect 537254 565214 543322 567414
rect 510541 565014 510542 565214
rect 510742 565014 543322 565214
rect 510541 565013 510743 565014
rect 327239 560030 327441 560031
rect 297340 559830 327240 560030
rect 327440 559830 327441 560030
rect 297340 557630 303408 559830
rect 327239 559829 327441 559830
rect 510631 560030 510833 560031
rect 537254 560030 543322 565014
rect 510631 559830 510632 560030
rect 510832 559830 543322 560030
rect 510631 559829 510833 559830
rect 327233 557630 327435 557631
rect 297340 557430 327234 557630
rect 327434 557430 327435 557630
rect 297340 555230 303408 557430
rect 327233 557429 327435 557430
rect 510645 557630 510847 557631
rect 537254 557630 543322 559830
rect 510645 557430 510646 557630
rect 510846 557430 543322 557630
rect 510645 557429 510847 557430
rect 327233 555230 327435 555231
rect 297340 555030 327234 555230
rect 327434 555030 327435 555230
rect 297340 552830 303408 555030
rect 327233 555029 327435 555030
rect 510627 555230 510829 555231
rect 537254 555230 543322 557430
rect 510627 555030 510628 555230
rect 510828 555030 543322 555230
rect 510627 555029 510829 555030
rect 327237 552830 327439 552831
rect 297340 552630 327238 552830
rect 327438 552630 327439 552830
rect 297340 550430 303408 552630
rect 327237 552629 327439 552630
rect 510623 552830 510825 552831
rect 537254 552830 543322 555030
rect 510623 552630 510624 552830
rect 510824 552630 543322 552830
rect 510623 552629 510825 552630
rect 327217 550430 327419 550431
rect 297340 550230 327218 550430
rect 327418 550230 327419 550430
rect 297340 548030 303408 550230
rect 327217 550229 327419 550230
rect 510617 550430 510819 550431
rect 537254 550430 543322 552630
rect 510617 550230 510618 550430
rect 510818 550230 543322 550430
rect 510617 550229 510819 550230
rect 327219 548030 327421 548031
rect 297340 547830 327220 548030
rect 327420 547830 327421 548030
rect 297340 515792 303408 547830
rect 327219 547829 327421 547830
rect 510605 548030 510807 548031
rect 537254 548030 543322 550230
rect 510605 547830 510606 548030
rect 510806 547830 543322 548030
rect 510605 547829 510807 547830
rect 537254 515792 543322 547830
rect 297218 509724 543322 515792
<< via4 >>
rect 578435 644584 580895 644585
rect 569603 642244 572065 642245
rect 569603 639784 569604 642244
rect 569604 639784 572064 642244
rect 572064 639784 572065 642244
rect 578435 642124 578436 644584
rect 578436 642124 580895 644584
rect 578435 642123 580895 642124
rect 569603 639783 572065 639784
rect 572603 634584 575063 634585
rect 572603 632124 572604 634584
rect 572604 632124 575063 634584
rect 572603 632123 575063 632124
rect 576893 632244 579353 632245
rect 576893 629784 576894 632244
rect 576894 629784 579353 632244
rect 576893 629783 579353 629784
rect 327364 598348 327716 598700
rect 516340 598224 516692 598576
rect 327836 595038 328188 595390
rect 510484 595038 510836 595390
rect 327716 591038 328068 591390
rect 510446 591038 510798 591390
rect 327368 587038 327720 587390
rect 511122 587038 511474 587390
rect 327878 583038 328230 583390
rect 510472 583038 510824 583390
rect 510464 579038 510816 579390
rect 327506 578338 327858 578690
rect 327464 575038 327816 575390
rect 510510 575038 510862 575390
rect 327534 571038 327886 571390
rect 510456 571038 510808 571390
rect 326860 566776 327212 567128
rect 510918 566754 511270 567106
<< metal5 >>
rect 287400 597414 293468 650884
rect 546148 644584 552216 650962
rect 578411 644585 580919 644609
rect 578411 644584 578435 644585
rect 546148 642245 578435 644584
rect 546148 639784 569603 642245
rect 546148 634584 552216 639784
rect 569579 639783 569603 639784
rect 572065 642124 578435 642245
rect 572065 639783 572089 642124
rect 578411 642123 578435 642124
rect 580895 642123 580919 644585
rect 578411 642099 580919 642123
rect 569579 639759 572089 639783
rect 572579 634585 575087 634609
rect 572579 634584 572603 634585
rect 546148 632123 572603 634584
rect 575063 632244 575087 634585
rect 576869 632245 579377 632269
rect 576869 632244 576893 632245
rect 575063 632123 576893 632244
rect 546148 629784 576893 632123
rect 327340 599014 329382 599414
rect 509068 599014 516716 599414
rect 327340 598700 327740 599014
rect 327340 598348 327364 598700
rect 327716 598348 327740 598700
rect 327340 598324 327740 598348
rect 516316 598576 516716 599014
rect 516316 598224 516340 598576
rect 516692 598224 516716 598576
rect 516316 598200 516716 598224
rect 546148 597414 552216 629784
rect 576869 629783 576893 629784
rect 579353 629783 579377 632245
rect 576869 629759 579377 629783
rect 287400 597014 329382 597414
rect 509068 597014 552216 597414
rect 287400 593414 293468 597014
rect 327812 595390 329382 595414
rect 327812 595038 327836 595390
rect 328188 595038 329382 595390
rect 327812 595014 329382 595038
rect 509068 595390 510860 595414
rect 509068 595038 510484 595390
rect 510836 595038 510860 595390
rect 509068 595014 510860 595038
rect 546148 593414 552216 597014
rect 287400 593014 329382 593414
rect 509068 593014 552216 593414
rect 287400 589414 293468 593014
rect 327692 591390 329382 591414
rect 327692 591038 327716 591390
rect 328068 591038 329382 591390
rect 327692 591014 329382 591038
rect 509068 591390 510822 591414
rect 509068 591038 510446 591390
rect 510798 591038 510822 591390
rect 509068 591014 510822 591038
rect 546148 589414 552216 593014
rect 287400 589014 329382 589414
rect 509068 589014 552216 589414
rect 287400 585414 293468 589014
rect 327344 587390 329382 587414
rect 327344 587038 327368 587390
rect 327720 587038 329382 587390
rect 327344 587014 329382 587038
rect 509068 587390 511498 587414
rect 509068 587038 511122 587390
rect 511474 587038 511498 587390
rect 509068 587014 511498 587038
rect 546148 585414 552216 589014
rect 287400 585014 329382 585414
rect 509068 585014 552216 585414
rect 287400 581414 293468 585014
rect 327854 583390 329382 583414
rect 327854 583038 327878 583390
rect 328230 583038 329382 583390
rect 327854 583014 329382 583038
rect 509068 583390 510848 583414
rect 509068 583038 510472 583390
rect 510824 583038 510848 583390
rect 509068 583014 510848 583038
rect 546148 581414 552216 585014
rect 287400 581014 329382 581414
rect 509068 581014 552216 581414
rect 287400 577414 293468 581014
rect 327482 579014 329382 579414
rect 509068 579390 510840 579414
rect 509068 579038 510464 579390
rect 510816 579038 510840 579390
rect 509068 579014 510840 579038
rect 327482 578690 327882 579014
rect 327482 578338 327506 578690
rect 327858 578338 327882 578690
rect 327482 578314 327882 578338
rect 546148 577414 552216 581014
rect 287400 577014 329382 577414
rect 509068 577014 552216 577414
rect 287400 573414 293468 577014
rect 327440 575390 329382 575414
rect 327440 575038 327464 575390
rect 327816 575038 329382 575390
rect 327440 575014 329382 575038
rect 509068 575390 510886 575414
rect 509068 575038 510510 575390
rect 510862 575038 510886 575390
rect 509068 575014 510886 575038
rect 546148 573414 552216 577014
rect 287400 573014 329382 573414
rect 509068 573014 552216 573414
rect 287400 569414 293468 573014
rect 327510 571390 329382 571414
rect 327510 571038 327534 571390
rect 327886 571038 329382 571390
rect 327510 571014 329382 571038
rect 509068 571390 510832 571414
rect 509068 571038 510456 571390
rect 510808 571038 510832 571390
rect 509068 571014 510832 571038
rect 546148 569414 552216 573014
rect 287400 569014 329382 569414
rect 509068 569014 552216 569414
rect 287400 565414 293468 569014
rect 326836 567128 329382 567414
rect 326836 566776 326860 567128
rect 327212 567014 329382 567128
rect 509068 567106 511294 567414
rect 509068 567014 510918 567106
rect 327212 566776 327236 567014
rect 326836 566752 327236 566776
rect 510894 566754 510918 567014
rect 511270 566754 511294 567106
rect 510894 566730 511294 566754
rect 546148 565414 552216 569014
rect 287400 565014 329382 565414
rect 509068 565014 552216 565414
rect 287400 504794 293468 565014
rect 546148 504794 552216 565014
rect 287400 498726 552216 504794
rect 287400 498714 293468 498726
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
<< end >>
